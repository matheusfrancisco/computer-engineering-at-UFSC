*Netlist_teste
Vgs1 in N001 AC 1 
VGS N001 0 1.2067 
M§N_1u Vout in 0 0 N_1u l=4.0697u w=63.2713u 
RD VDD Vout 40688.4657 
VDS VDD 0 5V 
.model NMOS NMOS 
.model PMOS PMOS 
.lib C:\Program Files (x86)\LTC\LTspiceIV\lib\cmp\standard.mos 
.include cmosedu_models.txt 
.ac dec 10 1 1Mega
.measure AC GAIN FIND V(vout) AT = 1 
.backanno 
.end 
