*Netlist_teste
Vgs1 in N001 AC 1 
VGS N001 0 4.4572 
M§N_1u Vout in 0 0 N_1u l=4.5676u w=9.7645u 
RD VDD Vout 10868.1317 
VDS VDD 0 5V 
.model NMOS NMOS 
.model PMOS PMOS 
.lib C:\Program Files (x86)\LTC\LTspiceIV\lib\cmp\standard.mos 
.include cmosedu_models.txt 
.ac dec 10 1 1Mega
.measure AC GAIN FIND V(vout) AT = 1 
.backanno 
.end 
