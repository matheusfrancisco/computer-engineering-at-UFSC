*Netlist_teste
Vd Vdd 0 5V 
M1 Vdd N001 N001 Vdd P_1u l=20.000000u w=3.000000u 
M2 Vdd N001 vout Vdd P_1u l=20.000000u w=3.000000u 
Iref N001 0 137812.297564uA
M3 vout N002 0 0 N_1u l=1.500000u w=3.000000u 
VGS N003 0 1.363323
Vg N002 N003 AC 1
.model NMOS NMOS
.model PMOS PMOS
.lib C:\Program Files (x86)\LTC\LTspiceIV\lib\cmp\standard.mos
.ac oct 1 1 1MEG
.include cmosedu_models.txt 
.meas AC gain FIND V(vout) AT 1 
.backanno 
.end 
