
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_SIGNED.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;


entity ROM is
Generic (
	      --
		   -- Size of the address bus.
		   --
		   p_ROM_SIZE		 : integer := 4				
	 );
    Port ( 
				i_CLK			 : in STD_LOGIC;
				i_EN 			 : in STD_LOGIC;
				i_ADDRESS    : in STD_LOGIC_VECTOR ((p_ROM_SIZE-1) downto 0);
				o_DATA       : out STD_LOGIC_VECTOR (31 downto 0));
end ROM;

architecture Behavioral of ROM is
-------------------------------------------------------------------------------------
-- Sinais internos e componentes.
-------------------------------------------------------------------------------------
--	signal i : integer;
	
	type ROM_TYPE is array(0 TO ((2**p_ROM_SIZE)-1)) of std_logic_vector(o_DATA'range);
 
    signal ROM : ROM_TYPE := (
    x"50000003", -- 0101 0010 0000 0000 0000 0000 0000 0011
    x"52000002", 
    x"1E200000", -- 0001 1110 0010 0000 0000 0000 0000 0000
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000",
	 
	 x"00000000", -- 0101 0010 0000 0000 0000 0000 0000 0011
    x"00000000", 
    x"00000000", -- 0001 1110 0010 0000 0000 0000 0000 0000
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000",

    x"00000000", -- 0101 0010 0000 0000 0000 0000 0000 0011
    x"00000000", 
    x"00000000", -- 0001 1110 0010 0000 0000 0000 0000 0000
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000",

    x"00000000", -- 0101 0010 0000 0000 0000 0000 0000 0011
    x"00000000", 
    x"00000000", -- 0001 1110 0010 0000 0000 0000 0000 0000
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000", 
    x"00000000"	 
    );
 
    attribute rom_style : string;
    attribute rom_style of ROM : signal is "block"; 
  
-------------------------------------------------------------------------------------
begin
-------------------------------------------------------------------------------------

	PROCESS(i_CLK)
	BEGIN
		IF RISING_EDGE(i_CLK) THEN
			IF (i_EN = '1') THEN
				o_DATA <= ROM(conv_integer(i_ADDRESS));
			END IF;
		END IF;
	END PROCESS;

end Behavioral;